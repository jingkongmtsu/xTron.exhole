Coord:     0.000000      0.000000      5.272336
Rho  GAA  TA  LA
    0.00000005923267     0.00000000000004     0.00000015901972     0.00000060713751
    0.37500000000000     -0.00000007473237
    6.00000000000000     -0.00061963376273
Coord:     0.000000      0.000000      0.065091
Rho  GAA  TA  LA
    1.39121591611408    25.72901643566057     4.62347651030445  -179.27936980288987
    0.37500000000000     -0.42421026580810
    6.00000000000000     -0.00000000674660
Coord:     0.000000      0.000000      0.585815
Rho  GAA  TA  LA
    0.20154948535548     0.48780817303610     0.60507246170306     0.03584309073940
    0.37500000000000     -0.20035545546576
    6.00000000000000     -0.00000000998692
